/*
    нс - наносекунди
    мс - мілісекунди
    СІ - семисегментний індикатор

    В цьому файлі проведу симуляцію свого модуля, що керує СІ.
    Цей модуль тактується частотою 50 МГц і керує чотирьма СІ.

    За однин період він почергово драйвить всі 4 СІ. Період його роботи це 50 000 тактів, ...
    на частоті в 50 МГц це 10 мс. Таким чином кожен СІ драйвиться 2,5 мс, а чстота драйву ...
    складає 100 Гц. Для сприйняття людиною цього достатньо. 

    Буду симулювати протягом однієї секунди. На цьому проміжку буде два ресети.



*/


// Встановлюю частові координати
`timescale 1ns/100ps

module tb_for_selector ();

    reg clk_i = 0;
    reg rst_n_i;
    reg [15:0] reg_16_i;
    wire [6:0] seg_display_o;
    wire [3:0] SS_o;


    parameter P = 20;   // Період становить 20 нс, тобто частота 50 МГц
    parameter Tms = P * 50 * 1000; // Часовий проміжок в одну мс

    // Екземпляр модуля декодера
    selector selector_inst(
        .clk_i(clk_i),
        .rst_n_i(rst_n_i),
        .reg_16_i(reg_16_i),
        .seg_display_o(seg_display_o),
        .SS_o(SS_o)
    );


    initial # (Tms * 100) $stop; // Моделювання триватиме 100мс


    initial forever #(P / 2) clk_i = ~clk_i; // Формую тактовий сигнал


    // Гереування ресетів
    initial begin
        // Перший ресет на 10мс від початку симуляції. 
        # (Tms * 10)
        # (Tms) rst_n_i = 1;
        # (Tms) rst_n_i = 0;
        # (Tms) rst_n_i = 1;

        // Тут вже пройшло 13 мс. Другий ресет на 60 мс
        # (Tms * 47)
        # (Tms) rst_n_i = 1;
        # (Tms) rst_n_i = 0;
        # (Tms) rst_n_i = 1;
    end

    // Гереування інформації для СІ
    initial begin  
        // На 20 мс
        # (Tms * 20)
        reg_16_i = 16'b0;

        // На 40мс
        # (Tms * 20)
        reg_16_i = 16'h1234;

        // На 60мс
        # (Tms * 20)
        reg_16_i = 16'h4321;

         // На 80мс
        # (Tms * 20)
        reg_16_i = 16'hFEDC;
    end
    
endmodule
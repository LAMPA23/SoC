
module ES (
	clk_clk,
	reset_reset_n,
	to_leds_readdata);	

	input		clk_clk;
	input		reset_reset_n;
	output	[31:0]	to_leds_readdata;
endmodule
